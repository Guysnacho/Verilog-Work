module top(A, B, C, D, F);

input A, B, C, D;
output F;

// YOUR VERILOG CODE BELOW

endmodule
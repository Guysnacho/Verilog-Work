// starter.v (Rename to <RNumber>.v
//
// Implement an 32-to-1 Decoder
//
module top(S, I, Y)

// Verilog Code Here.

endmodule

// Additional Modules Here (if needed).
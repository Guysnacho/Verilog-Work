// starter.v (RENAME TO <RNumber>.v
//
// Implement a 5-to-32 Line Decoder.
//

module top(A, D)

// YOUR VERILOG CODE HERE

endmodule

// OTHER MODULES HERE (IF REQUIRED)
// starter.v (Rename to <RNumber>.v
//
//  Implement an 8-bit Adder Subtractor.
//
module top(Cin, A, B, Cout, S)

// Verilog code goes here.

endmodule

// Additional modules go here (if necessary).